library verilog;
use verilog.vl_types.all;
entity Control_Unit_tb is
end Control_Unit_tb;
