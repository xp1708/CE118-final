library verilog;
use verilog.vl_types.all;
entity RegisterFile_vlg_vec_tst is
end RegisterFile_vlg_vec_tst;
