library verilog;
use verilog.vl_types.all;
entity giaithua_vlg_vec_tst is
end giaithua_vlg_vec_tst;
