library verilog;
use verilog.vl_types.all;
entity One_Counter_tb is
end One_Counter_tb;
