library verilog;
use verilog.vl_types.all;
entity mux16_1_vlg_vec_tst is
end mux16_1_vlg_vec_tst;
