library verilog;
use verilog.vl_types.all;
entity Data_Path_vlg_vec_tst is
end Data_Path_vlg_vec_tst;
