module comp(a,comp);
	input wire [15:0] a;
	output [15:0]comp; 
	assign comp = a;
endmodule