library verilog;
use verilog.vl_types.all;
entity Lab01_CE118_22521154_vlg_check_tst is
    port(
        LEDG1           : in     vl_logic;
        LEDG2           : in     vl_logic;
        LEGG0           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab01_CE118_22521154_vlg_check_tst;
