library verilog;
use verilog.vl_types.all;
entity parallel_datapath_vlg_vec_tst is
end parallel_datapath_vlg_vec_tst;
