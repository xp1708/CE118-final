library verilog;
use verilog.vl_types.all;
entity controler_vlg_vec_tst is
end controler_vlg_vec_tst;
