library verilog;
use verilog.vl_types.all;
entity RF_vlg_vec_tst is
end RF_vlg_vec_tst;
