library verilog;
use verilog.vl_types.all;
entity Moore_Detector_vlg_vec_tst is
end Moore_Detector_vlg_vec_tst;
