library verilog;
use verilog.vl_types.all;
entity Counter_tb is
end Counter_tb;
