library verilog;
use verilog.vl_types.all;
entity Lab01_CE118_22521154 is
    port(
        LEDG2           : out    vl_logic;
        SW2             : in     vl_logic;
        KEY1            : in     vl_logic;
        SW0             : in     vl_logic;
        SW1             : in     vl_logic;
        KEY0            : in     vl_logic;
        LEDG1           : out    vl_logic;
        LEGG0           : out    vl_logic
    );
end Lab01_CE118_22521154;
