library verilog;
use verilog.vl_types.all;
entity Top_module_vlg_vec_tst is
end Top_module_vlg_vec_tst;
