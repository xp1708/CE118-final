library verilog;
use verilog.vl_types.all;
entity Lab01_CE118_22521154_vlg_vec_tst is
end Lab01_CE118_22521154_vlg_vec_tst;
