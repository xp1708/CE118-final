library verilog;
use verilog.vl_types.all;
entity Data_Path is
    port(
        CLK             : in     vl_logic;
        DataIn          : in     vl_logic_vector(15 downto 0);
        IE              : in     vl_logic;
        WAA             : in     vl_logic_vector(3 downto 0);
        WEA             : in     vl_logic;
        WAB             : in     vl_logic_vector(3 downto 0);
        WEB             : in     vl_logic;
        RAA             : in     vl_logic_vector(3 downto 0);
        REA             : in     vl_logic;
        RAB             : in     vl_logic_vector(3 downto 0);
        REB             : in     vl_logic;
        OE              : in     vl_logic;
        S_ALU1          : in     vl_logic_vector(3 downto 0);
        S_ALU2          : in     vl_logic_vector(3 downto 0);
        \Out\           : out    vl_logic_vector(15 downto 0);
        Datapath        : out    vl_logic_vector(15 downto 0);
        mux_to_rf       : out    vl_logic_vector(15 downto 0)
    );
end Data_Path;
