module mux2_1(a,b,sel,muxout);
	input [15:0]a;
	input [15:0]b;
	input sel;
	output [15:0]muxout;
	
	assign muxout = (sel) ? a: b;
endmodule