my_counter_inst : my_counter PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
