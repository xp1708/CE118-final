library verilog;
use verilog.vl_types.all;
entity shiftleft_vlg_vec_tst is
end shiftleft_vlg_vec_tst;
