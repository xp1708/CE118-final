library verilog;
use verilog.vl_types.all;
entity One_Counter_vlg_vec_tst is
end One_Counter_vlg_vec_tst;
