module FullAdder(a,b,ci,s,add_overflow,zero);
	input wire [3:0] a;
	input wire [3:0] b;
	input wire ci;
	wire co0, co1, co2, co3;
	output wire [3:0] s;
	output wire add_overflow;
	output wire zero;
	
	assign co0 = (ci&a[0]) | (ci&b[0]) | (a[0]&b[0]);
	assign s[0] = a[0]^b[0]^ci;
	
	assign co1 = (co0&a[1]) | (co0&b[1]) | (a[1]&b[1]);
	assign s[1] = a[1]^b[1]^co0;
	
	assign co2 = (co1&a[2]) | (co1&b[2]) | (a[2]&b[2]);
	assign s[2] = a[2]^b[2]^co1;
	
	assign co3 = (co2&a[3]) | (co2&b[3]) | (a[3]&b[3]);
	assign s[3] = a[3]^b[3]^co2;
	
	assign add_overflow = (co2 ^ co3);
	assign zero = (s==4'b0000);
	
	
endmodule