library verilog;
use verilog.vl_types.all;
entity detector_Mealy_vlg_vec_tst is
end detector_Mealy_vlg_vec_tst;
