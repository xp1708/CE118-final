library verilog;
use verilog.vl_types.all;
entity detector_vlg_vec_tst is
end detector_vlg_vec_tst;
