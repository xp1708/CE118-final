library verilog;
use verilog.vl_types.all;
entity one_counter_op_vlg_vec_tst is
end one_counter_op_vlg_vec_tst;
