library verilog;
use verilog.vl_types.all;
entity Lab01_CE118_22521154_vlg_sample_tst is
    port(
        KEY0            : in     vl_logic;
        KEY1            : in     vl_logic;
        SW0             : in     vl_logic;
        SW1             : in     vl_logic;
        SW2             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Lab01_CE118_22521154_vlg_sample_tst;
