module comp(a,comp);
	input wire [3:0] a;
	output [3:0]comp; 
	assign comp = a;
endmodule